library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cpu_test is
end cpu_test;

architecture cpu_test of cpu_test is
begin
end cpu_test;
